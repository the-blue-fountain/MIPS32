`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.09.2024 12:53:25
// Design Name: 
// Module Name: left_shift_32bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module left_shift_32bit(out,a,b);
    input [31:0] a;
    input [4:0] b;
    output [31:0] out;
    wire [31:0] t[31:0];

    assign t[0]={31'b0,a[0]};
    assign t[1]={30'b0,a[0],a[1]};
    assign t[2]={29'b0,a[0],a[1],a[2]};
    assign t[3]={28'b0,a[0],a[1],a[2],a[3]};
    assign t[4]={27'b0,a[0],a[1],a[2],a[3],a[4]};
    assign t[5]={26'b0,a[0],a[1],a[2],a[3],a[4],a[5]};
    assign t[6]={25'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6]};
    assign t[7]={24'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7]};
    assign t[8]={23'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8]};
    assign t[9]={22'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9]};
    assign t[10]={21'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10]};
    assign t[11]={20'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11]};
    assign t[12]={19'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12]};
    assign t[13]={18'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13]};
    assign t[14]={17'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14]};
    assign t[15]={16'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15]};
    assign t[16]={15'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16]};
    assign t[17]={14'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17]};
    assign t[18]={13'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18]};
    assign t[19]={12'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19]};
    assign t[20]={11'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20]};
    assign t[21]={10'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21]};
    assign t[22]={9'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22]};
    assign t[23]={8'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23]};
    assign t[24]={7'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24]};
    assign t[25]={6'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25]};
    assign t[26]={5'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25],a[26]};
    assign t[27]={4'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25],a[26],a[27]};
    assign t[28]={3'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25],a[26],a[27],a[28]};
    assign t[29]={2'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25],a[26],a[27],a[28],a[29]};
    assign t[30]={1'b0,a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25],a[26],a[27],a[28],a[29],a[30]};
    assign t[31]={a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[16],a[17],a[18],a[19],a[20],a[21],a[22],a[23],a[24],a[25],a[26],a[27],a[28],a[29],a[30],a[31]};
    
    MUX_32_to_1 M0(out[0],b,t[0]);
    MUX_32_to_1 M1(out[1],b,t[1]);
    MUX_32_to_1 M2(out[2],b,t[2]);
    MUX_32_to_1 M3(out[3],b,t[3]);
    MUX_32_to_1 M4(out[4],b,t[4]);
    MUX_32_to_1 M5(out[5],b,t[5]);
    MUX_32_to_1 M6(out[6],b,t[6]);
    MUX_32_to_1 M7(out[7],b,t[7]);
    MUX_32_to_1 M8(out[8],b,t[8]);
    MUX_32_to_1 M9(out[9],b,t[9]);
    MUX_32_to_1 M10(out[10],b,t[10]);
    MUX_32_to_1 M11(out[11],b,t[11]);
    MUX_32_to_1 M12(out[12],b,t[12]);
    MUX_32_to_1 M13(out[13],b,t[13]);
    MUX_32_to_1 M14(out[14],b,t[14]);
    MUX_32_to_1 M15(out[15],b,t[15]);
    MUX_32_to_1 M16(out[16],b,t[16]);
    MUX_32_to_1 M17(out[17],b,t[17]);
    MUX_32_to_1 M18(out[18],b,t[18]);
    MUX_32_to_1 M19(out[19],b,t[19]);
    MUX_32_to_1 M20(out[20],b,t[20]);
    MUX_32_to_1 M21(out[21],b,t[21]);
    MUX_32_to_1 M22(out[22],b,t[22]);
    MUX_32_to_1 M23(out[23],b,t[23]);
    MUX_32_to_1 M24(out[24],b,t[24]);
    MUX_32_to_1 M25(out[25],b,t[25]);
    MUX_32_to_1 M26(out[26],b,t[26]);
    MUX_32_to_1 M27(out[27],b,t[27]);
    MUX_32_to_1 M28(out[28],b,t[28]);
    MUX_32_to_1 M29(out[29],b,t[29]);
    MUX_32_to_1 M30(out[30],b,t[30]);
    MUX_32_to_1 M31(out[31],b,t[31]);
endmodule
